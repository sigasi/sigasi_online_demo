------------------------------------------------------------------------------------------------------------------------
-- If you got this far, you have learned the basics about working with Sigasi Studio for VS Code.
--
-- Congratulations!
--
-- You are now ready to go and set up a project for your own VHDL code.
------------------------------------------------------------------------------------------------------------------------
-- If you were to encounter any issues you can contact us at support@sigasi.com
--
-- You can find the Sigasi logs by opening the log and tracing log view.
-- Open the `Command Palette (Ctrl+Shift+P)` and type `Sigasi: Open log` or `Sigasi: Open log`.
--
-- To increase the logging in the Sigasi log view you can increase the level of logging the server produces
-- by opening the `Command Palette (Ctrl+Shift+P)` and typing `Sigasi: Set the log level of the Sigasi language server`.
-- `info` is usually enough information for us.
--
-- To see all the tracing logs you should open the settings and set `Sigasi>trace:server` to `verbose`.
------------------------------------------------------------------------------------------------------------------------



------------------------------------------------------------------------------------------------------------------------
-- NEXT STEPS
--
-- Now browse folders tb, vhdl and vlog and open the design files in those folders.
-- Note that tb folder has the file testbench.sv which instatiates a module named cmd_gen.
-- Also view the components that are instatiated by cmd_gen module and go through the TODOs in those design files.
------------------------------------------------------------------------------------------------------------------------